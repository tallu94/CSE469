// EE469 LAB 1
// Erika Burk, Jeff Josephsen, Ameer Talal Mahmood

module instruction_decoder (instruction_set, rm, shift, rn, rd, rotate, immediateValue,
		 br_address, dt_address, ALUCtl_code, enable, execute_flag );

	input wire  [31:0] instruction_set;
	input wire enable;

	output wire [3:0]  rm;
	output wire [7:0]  shift;
	output wire [3:0]  rn;
	output wire [3:0]  rd;
	output wire [3:0]	rotate;					// shift applied to an immediate value
	output wire [7:0]  immediateValue;
	wire [3:0]  cond_field;				// flags for alu
	output wire [23:0] br_address;				// address to branch 
	output wire [11:0] dt_address;  			// used in LDR and STR as an immediate offset
	output wire [10:0] ALUCtl_code;

	input wire [31:0] cpsr;
	output wire execute_flag; 					//if condition field matches cpsr, true, else false

	assign cond_field = instruction_set[31:28];

/* 	initial begin
		rm = 4'b0;
		shift = 11'b0;
		rn = 4'b0;
		rd = 4'b0;
		immediateValue = 8'b0;
		dt_address = 12'b0;
		br_address = 24'bx;
		cond_field = 4'b0;
		ALUCtl_code = 11'dx;		// initial ALU state (does nothing)
	end */

	// case statememt to decode instruction set
	always @(*) begin

		if (enable) begin

			case (cond_field)
				4'b0000: execute_flag = cpsr[30];
				4'b0001: execute_flag = ~cpsr[30];
				4'b0010: execute_flag = cpsr[29];
				4'b0011: execute_flag = ~cpsr[29];
				4'b0100: execute_flag = cpsr[31];
				4'b0101: execute_flag = ~cpsr[31];
				4'b0110: execute_flag = cpsr[28];
				4'b0111: execute_flag = ~cpsr[28];
				4'b1000: execute_flag = cpsr[29] & ~cpsr[30];
				4'b1001: execute_flag = ~cpsr[29] & cpsr[30];
				4'b1010: execute_flag = (cpsr[31] & cpsr[28]) | (~cpsr[31] & ~cpsr[28]); 
				4'b1011: execute_flag = (cpsr[31] & ~cpsr[28]) | (~cpsr[31] & cpsr[28]);
				4'b1100: execute_flag = ~cpsr[30] & ((cpsr[31] & cpsr[28]) | (~cpsr[31] & ~cpsr[28]));
				4'b1101: execute_flag = cpsr[30] | (cpsr[31] & ~cpsr[28]) | (~cpsr[31] & cpsr[28]);
				4'b1110: execute_flag = 1'b1;
				default: execute_flag = 1'b1;
			endcase

			casex(instruction_set[27:20])

				// ------------- DATA PROCESSING OPERATIONS (0-30) --------------
				8'b0000100x: begin 						// ADD
					rm = instruction_set[3:0];
					shift = instruction_set[11:4];
					rn = instruction_set[19:16];
					rd = instruction_set[15:12];
					rotate = 4'bx;
					immediateValue = 8'bx;
					dt_address = 12'bx;
					br_address = 24'bx;
					cond_field = instruction_set[31:28];
					ALUCtl_code = 11'd0;
				end

				8'b0010100x: begin 						// ADDI
					rm = 4'bx;
					shift = instruction_set[11:4];
					rn = instruction_set[19:16];
					rd = instruction_set[15:12];
					rotate = 4'bx;
					immediateValue = instruction_set[7:0];
					dt_address = 12'bx;
					br_address = 24'bx;
					cond_field = instruction_set[31:28];
					ALUCtl_code = 11'd1;
				end

				8'b0000010x: begin 						// SUB
					rm = instruction_set[3:0];
					shift = instruction_set[11:4];
					rn = instruction_set[19:16];
					rd = instruction_set[15:12];
					rotate = 4'bx;
					immediateValue = 8'bx;
					dt_address = 12'bx;
					br_address = 24'bx;
					cond_field = instruction_set[31:28];
					ALUCtl_code = 11'd2;
				end

				8'b0000000x: begin 						// AND
					rm = instruction_set[3:0];
					shift = instruction_set[11:4];
					rn = instruction_set[19:16];
					rd = instruction_set[15:12];
					rotate = 4'bx;
					immediateValue = 8'bx;
					dt_address = 12'bx;
					br_address = 24'bx;
					cond_field = instruction_set[31:28];
					ALUCtl_code = 11'd3;
				end

				8'b0001100x: begin 						// ORR
					rm = instruction_set[3:0];
					shift = instruction_set[11:4];
					rn = instruction_set[19:16];
					rd = instruction_set[15:12];
					rotate = 4'bx;
					immediateValue = 8'bx;
					dt_address = 12'bx;
					br_address = 24'bx;
					cond_field = instruction_set[31:28];
					ALUCtl_code = 11'd4;
				end

				8'b0000001x: begin 						// EOR
					rm = instruction_set[3:0];
					shift = instruction_set[11:4];
					rn = instruction_set[19:16];
					rd = instruction_set[15:12];
					rotate = 4'bx;
					immediateValue = 8'bx;
					dt_address = 12'bx;
					br_address = 24'bx;
					cond_field = instruction_set[31:28];
					ALUCtl_code = 11'd5;
				end

				8'b0001101x: begin 						// MOV
					rm = instruction_set[3:0];
					shift = instruction_set[11:4];
					rn = instruction_set[19:16];
					rd = instruction_set[15:12];
					rotate = 4'bx;
					immediateValue = 8'bx;
					dt_address = 12'bx;
					br_address = 24'bx;
					cond_field = instruction_set[31:28];
					ALUCtl_code = 11'd6;
				end

				8'b0001111x: begin 						// MNV
					rm = instruction_set[3:0];
					shift = instruction_set[11:4];
					rn = instruction_set[19:16];
					rd = instruction_set[15:12];
					rotate = 4'bx;
					immediateValue = 8'bx;
					dt_address = 12'bx;
					br_address = 24'bx;
					cond_field = instruction_set[31:28];
					ALUCtl_code = 11'd7;
				end

				8'b0001010x: begin 						// CMP
					rm = instruction_set[3:0];
					shift = instruction_set[11:4];
					rn = instruction_set[19:16];
					rd = instruction_set[15:12];
					rotate = 4'bx;
					immediateValue = 8'bx;
					dt_address = 12'bx;
					br_address = 24'bx;
					cond_field = instruction_set[31:28];
					ALUCtl_code = 11'd8;
				end

				8'b0001000x: begin 						// TST
					rm = instruction_set[3:0];
					shift = instruction_set[11:4];
					rn = instruction_set[19:16];
					rd = instruction_set[15:12];
					rotate = 4'bx;
					immediateValue = 8'bx;
					dt_address = 12'bx;
					br_address = 24'bx;
					cond_field = instruction_set[31:28];
					ALUCtl_code = 11'd9;
				end

				8'b0001001x: begin 						// TEQ
					rm = instruction_set[3:0];
					shift = instruction_set[11:4];
					rn = instruction_set[19:16];
					rd = instruction_set[15:12];
					rotate = 4'bx;
					immediateValue = 8'bx;
					dt_address = 12'bx;
					br_address = 24'bx;
					cond_field = instruction_set[31:28];
					ALUCtl_code = 11'd10;
				end

				8'b0001110x: begin 						// BIC
					rm = instruction_set[3:0];
					shift = instruction_set[11:4];
					rn = instruction_set[19:16];
					rd = instruction_set[15:12];
					rotate = 4'bx;
					immediateValue = 8'bx;
					dt_address = 12'bx;
					br_address = 24'bx;
					cond_field = instruction_set[31:28];
					ALUCtl_code = 11'd11;
				end

				8'b0011101x: begin 						// MOVI
					rm = 4'bx;
					shift = 8'bx;
					rn = instruction_set[19:16];
					rd = instruction_set[15:12];
					rotate = instruction_set[11:8];
					immediateValue = instruction_set[7:0];
					dt_address = 12'bx;
					br_address = 24'bx;
					cond_field = instruction_set[31:28];
					ALUCtl_code = 11'd12;
				end

				8'b0011010x: begin 						// CMPI
					rm = 4'bx;
					shift = 8'bx;
					rn = instruction_set[19:16];
					rd = instruction_set[15:12];
					rotate = instruction_set[11:8];
					immediateValue = instruction_set[7:0];
					dt_address = 12'bx;
					br_address = 24'bx;
					cond_field = instruction_set[31:28];
					ALUCtl_code = 11'd13;
				end

				//------------- BRANCH/BRANCH-LINK (31-40) -----------------------
				8'b1010xxxx: begin 						// Branch
					rm = 4'bx;
					shift = 8'bx;
					rn = 4'bx;
					rd = 4'bx;
					rotate = 4'bx;
					immediateValue = 8'bx;
					dt_address = 12'bx;
					br_address = instruction_set[23:0];
					cond_field = instruction_set[31:28];
					ALUCtl_code = 11'd31;
				end

				8'b1011xxxx: begin 						// Branch and Link
					rm = 4'bx;
					shift = 8'bx;
					rn = 4'bx;
					rd = 4'bx;
					rotate = 4'bx;
					immediateValue = 8'bx;
					dt_address = 12'bx;
					br_address = instruction_set[23:0];
					cond_field = instruction_set[31:28];
					ALUCtl_code = 11'd32;				// use this later to determine when to BL in cpu.v to set R14
				end

				//------------- SINGLE DATA TRANSFER (41-50)----------------------
				8'b01xxxxx0: begin 						// LDR
					rm = instruction_set[3:0];
					shift = instruction_set[11:4];
					rn = instruction_set[19:16];
					rd = instruction_set[15:12];
					rotate = 4'bx;
					immediateValue = 8'bx;
					dt_address = instruction_set[23:0];
					br_address = 24'bx;
					cond_field = instruction_set[31:28];
					ALUCtl_code = 11'd41;
				end

				8'b01xxxxx1: begin 						// STR
					rm = instruction_set[3:0];
					shift = instruction_set[11:4];
					rn = instruction_set[19:16];
					rd = instruction_set[15:12];
					rotate = 4'bx;
					immediateValue = 8'bx;
					dt_address = instruction_set[23:0];
					br_address = 24'bx;
					cond_field = instruction_set[31:28];
					ALUCtl_code = 11'd42;
				end
				default: begin
					rm = 4'b0;
					shift = 11'b0;
					rn = 4'b0;
					rd = 4'b0;
					rotate = 4'bx;
					immediateValue = 8'b0;
					dt_address = 12'b0;
					br_address = 24'bx;
					cond_field = 4'b0;
					ALUCtl_code = 11'dx;
				end
			endcase
		end
	end
endmodule


/*module instruction_decoder_testbench();

	logic [31:0] instruction_set;
	logic [3:0]  rm;
	logic [7:0]  shift;
	logic [3:0]  rn;
	logic [3:0]  rd;
	logic [7:0] immediateValue;
	//output logic [3:0]	rotate;				// shift applied to an immediate value
	logic [3:0]  cond_field;				// flags for alu
	logic [23:0] br_address;				// address to branch to
	logic [11:0] dt_address;  			// used in LDR and STR as an immediate offset
	logic [10:0] ALUCtl_code;


  instruction_decoder dut(.instruction_set, .rm, .shift, .rn, .rd, .immediateValue, .cond_field,
			 .br_address, .dt_address, .ALUCtl_code);

  initial begin

  instruction_set =32'b11100000100001110101000000000110; #50	//ADD

	instruction_set =32'b11100001101000000000000000000011; #50 //MOV

	instruction_set =32'b11101010000000000000000000000000; #50 //b

	instruction_set =32'b11100010100001000100000000000001; #50	//ADDI

    $stop;

  end
endmodule*/