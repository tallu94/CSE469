library verilog;
use verilog.vl_types.all;
entity alu_testbench is
end alu_testbench;
