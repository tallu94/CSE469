library verilog;
use verilog.vl_types.all;
entity instruction_decoder_testbench is
end instruction_decoder_testbench;
