library verilog;
use verilog.vl_types.all;
entity test_testbench is
end test_testbench;
